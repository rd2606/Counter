`include "uvm_macros.svh"
import uvm_pkg::*;

`include "counter_transaction.sv"
`include "counter_sequencer.sv"
`include "counter_driver.sv"
`include "counter_monitor.sv"
`include "counter_agent.sv"
`include "counter_scoreboard.sv"
`include "counter_env.sv"
`include "counter_test.sv"
